module encoder_stateless (
	input signed [15:0] sample;
	input signed [15:0] 
);


	reg [15:0] step_sizes [89];
	wire [15:0] step;

	assign step = step_sizes[index];

endmodule
